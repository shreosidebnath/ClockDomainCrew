module EthMacDefinitions(
  input   clock,
  input   reset
);
endmodule
